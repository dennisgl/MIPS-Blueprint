library verilog;
use verilog.vl_types.all;
entity tb_SingleCycle is
end tb_SingleCycle;
